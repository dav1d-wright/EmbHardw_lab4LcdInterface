-- systemFile.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity systemFile is
	port (
		altpll_0_c2_clk            : out   std_logic;                                        --     altpll_0_c2.clk
		altpll_1_c0_clk            : out   std_logic;                                        --     altpll_1_c0.clk
		clk_clk                    : in    std_logic                     := '0';             --             clk.clk
		lcd_conduit_end_cs_n       : out   std_logic;                                        -- lcd_conduit_end.cs_n
		lcd_conduit_end_data       : inout std_logic_vector(15 downto 0) := (others => '0'); --                .data
		lcd_conduit_end_data_cmd_n : out   std_logic;                                        --                .data_cmd_n
		lcd_conduit_end_mode       : out   std_logic;                                        --                .mode
		lcd_conduit_end_rd_n       : out   std_logic;                                        --                .rd_n
		lcd_conduit_end_wr_n       : out   std_logic;                                        --                .wr_n
		lcd_conduit_end_lcdreset_n : out   std_logic;                                        --                .lcdreset_n
		reset_reset_n              : in    std_logic                     := '0';             --           reset.reset_n
		sdram_ctrl_wire_addr       : out   std_logic_vector(11 downto 0);                    -- sdram_ctrl_wire.addr
		sdram_ctrl_wire_ba         : out   std_logic_vector(1 downto 0);                     --                .ba
		sdram_ctrl_wire_cas_n      : out   std_logic;                                        --                .cas_n
		sdram_ctrl_wire_cke        : out   std_logic;                                        --                .cke
		sdram_ctrl_wire_cs_n       : out   std_logic;                                        --                .cs_n
		sdram_ctrl_wire_dq         : inout std_logic_vector(15 downto 0) := (others => '0'); --                .dq
		sdram_ctrl_wire_dqm        : out   std_logic_vector(1 downto 0);                     --                .dqm
		sdram_ctrl_wire_ras_n      : out   std_logic;                                        --                .ras_n
		sdram_ctrl_wire_we_n       : out   std_logic                                         --                .we_n
	);
end entity systemFile;

architecture rtl of systemFile is
	component systemFile_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(25 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			dtcm0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dtcm0_address                       : out std_logic_vector(25 downto 0);                    -- address
			dtcm0_read                          : out std_logic;                                        -- read
			dtcm0_clken                         : out std_logic;                                        -- clken
			dtcm0_write                         : out std_logic;                                        -- write
			dtcm0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			dtcm0_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			itcm0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			itcm0_address                       : out std_logic_vector(25 downto 0);                    -- address
			itcm0_read                          : out std_logic;                                        -- read
			itcm0_clken                         : out std_logic;                                        -- clken
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component systemFile_CPU;

	component LcdDriver is
		port (
			WaitReq_SO            : out   std_logic;                                        -- waitrequest
			Address_DI            : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			BurstCount_DI         : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			ByteEnable_DI         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			WriteData_DI          : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			ReadData_DO           : out   std_logic_vector(15 downto 0);                    -- readdata
			Read_SI               : in    std_logic                     := 'X';             -- read
			Write_SI              : in    std_logic                     := 'X';             -- write
			ReadDataValid_SO      : out   std_logic;                                        -- readdatavalid
			BeginBurstTransfer_SI : in    std_logic                     := 'X';             -- beginbursttransfer
			Clk_CI                : in    std_logic                     := 'X';             -- clk
			Reset_NRI             : in    std_logic                     := 'X';             -- reset_n
			Cs_NSO                : out   std_logic;                                        -- cs_n
			DB_DIO                : inout std_logic_vector(15 downto 0) := (others => 'X'); -- data
			DC_NSO                : out   std_logic;                                        -- data_cmd_n
			IM0_SO                : out   std_logic;                                        -- mode
			Rd_NSO                : out   std_logic;                                        -- rd_n
			Wr_NSO                : out   std_logic;                                        -- wr_n
			LcdReset_NRO          : out   std_logic                                         -- lcdreset_n
		);
	end component LcdDriver;

	component systemFile_SDRAM_ctrl is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(22 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component systemFile_SDRAM_ctrl;

	component systemFile_TCDM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component systemFile_TCDM;

	component systemFile_TCIM is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component systemFile_TCIM;

	component systemFile_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component systemFile_altpll_0;

	component systemFile_altpll_signalTap is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component systemFile_altpll_signalTap;

	component systemFile_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component systemFile_jtag_uart;

	component systemFile_performance_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component systemFile_performance_counter_0;

	component systemFile_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component systemFile_sysid;

	component systemFile_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component systemFile_timer_0;

	component systemFile_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                                    : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest                                : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                                       : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_readdatavalid                              : out std_logic;                                        -- readdatavalid
			CPU_data_master_write                                      : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address                             : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest                         : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read                                : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_master_readdatavalid                       : out std_logic;                                        -- readdatavalid
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			altpll_signalTap_pll_slave_address                         : out std_logic_vector(1 downto 0);                     -- address
			altpll_signalTap_pll_slave_write                           : out std_logic;                                        -- write
			altpll_signalTap_pll_slave_read                            : out std_logic;                                        -- read
			altpll_signalTap_pll_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_signalTap_pll_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_address                                : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                                  : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                                   : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess                            : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                          : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                           : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     : out std_logic;                                        -- chipselect
			LCD_avalon_slave_address                                   : out std_logic_vector(2 downto 0);                     -- address
			LCD_avalon_slave_write                                     : out std_logic;                                        -- write
			LCD_avalon_slave_read                                      : out std_logic;                                        -- read
			LCD_avalon_slave_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			LCD_avalon_slave_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			LCD_avalon_slave_beginbursttransfer                        : out std_logic;                                        -- beginbursttransfer
			LCD_avalon_slave_burstcount                                : out std_logic_vector(7 downto 0);                     -- burstcount
			LCD_avalon_slave_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			LCD_avalon_slave_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			LCD_avalon_slave_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			performance_counter_0_control_slave_address                : out std_logic_vector(4 downto 0);                     -- address
			performance_counter_0_control_slave_write                  : out std_logic;                                        -- write
			performance_counter_0_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_0_control_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_0_control_slave_begintransfer          : out std_logic;                                        -- begintransfer
			SDRAM_ctrl_s1_address                                      : out std_logic_vector(22 downto 0);                    -- address
			SDRAM_ctrl_s1_write                                        : out std_logic;                                        -- write
			SDRAM_ctrl_s1_read                                         : out std_logic;                                        -- read
			SDRAM_ctrl_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_ctrl_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_ctrl_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_ctrl_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_ctrl_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_ctrl_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sysid_control_slave_address                                : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TCIM_s2_address                                            : out std_logic_vector(9 downto 0);                     -- address
			TCIM_s2_write                                              : out std_logic;                                        -- write
			TCIM_s2_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TCIM_s2_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			TCIM_s2_byteenable                                         : out std_logic_vector(3 downto 0);                     -- byteenable
			TCIM_s2_chipselect                                         : out std_logic;                                        -- chipselect
			TCIM_s2_clken                                              : out std_logic;                                        -- clken
			timer_0_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                           : out std_logic;                                        -- write
			timer_0_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                      : out std_logic                                         -- chipselect
		);
	end component systemFile_mm_interconnect_0;

	component systemFile_mm_interconnect_1 is
		port (
			altpll_0_c0_clk                              : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			CPU_tightly_coupled_data_master_0_address    : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_tightly_coupled_data_master_0_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_tightly_coupled_data_master_0_read       : in  std_logic                     := 'X';             -- read
			CPU_tightly_coupled_data_master_0_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_tightly_coupled_data_master_0_write      : in  std_logic                     := 'X';             -- write
			CPU_tightly_coupled_data_master_0_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_tightly_coupled_data_master_0_clken      : in  std_logic                     := 'X';             -- clken
			TCDM_s1_address                              : out std_logic_vector(9 downto 0);                     -- address
			TCDM_s1_write                                : out std_logic;                                        -- write
			TCDM_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TCDM_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			TCDM_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			TCDM_s1_chipselect                           : out std_logic;                                        -- chipselect
			TCDM_s1_clken                                : out std_logic                                         -- clken
		);
	end component systemFile_mm_interconnect_1;

	component systemFile_mm_interconnect_2 is
		port (
			altpll_0_c0_clk                                   : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			CPU_tightly_coupled_instruction_master_0_address  : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_tightly_coupled_instruction_master_0_read     : in  std_logic                     := 'X';             -- read
			CPU_tightly_coupled_instruction_master_0_readdata : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_tightly_coupled_instruction_master_0_clken    : in  std_logic                     := 'X';             -- clken
			TCIM_s1_address                                   : out std_logic_vector(9 downto 0);                     -- address
			TCIM_s1_write                                     : out std_logic;                                        -- write
			TCIM_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TCIM_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			TCIM_s1_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			TCIM_s1_chipselect                                : out std_logic;                                        -- chipselect
			TCIM_s1_clken                                     : out std_logic                                         -- clken
		);
	end component systemFile_mm_interconnect_2;

	component systemFile_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component systemFile_irq_mapper;

	component systemfile_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component systemfile_rst_controller;

	component systemfile_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component systemfile_rst_controller_001;

	signal altpll_0_c0_clk                                                     : std_logic;                     -- altpll_0:c0 -> [CPU:clk, LCD:Clk_CI, SDRAM_ctrl:clk, TCDM:clk, TCIM:clk, TCIM:clk2, altpll_signalTap:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, mm_interconnect_2:altpll_0_c0_clk, performance_counter_0:clk, rst_controller:clk, sysid:clock, timer_0:clk]
	signal cpu_data_master_readdata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                         : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                         : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                             : std_logic_vector(25 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                          : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                                : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdatavalid                                       : std_logic;                     -- mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	signal cpu_data_master_write                                               : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                           : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                      : std_logic_vector(25 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                         : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata              : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest           : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                  : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                 : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_lcd_avalon_slave_beginbursttransfer               : std_logic;                     -- mm_interconnect_0:LCD_avalon_slave_beginbursttransfer -> LCD:BeginBurstTransfer_SI
	signal mm_interconnect_0_lcd_avalon_slave_readdata                         : std_logic_vector(15 downto 0); -- LCD:ReadData_DO -> mm_interconnect_0:LCD_avalon_slave_readdata
	signal mm_interconnect_0_lcd_avalon_slave_waitrequest                      : std_logic;                     -- LCD:WaitReq_SO -> mm_interconnect_0:LCD_avalon_slave_waitrequest
	signal mm_interconnect_0_lcd_avalon_slave_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:LCD_avalon_slave_address -> LCD:Address_DI
	signal mm_interconnect_0_lcd_avalon_slave_read                             : std_logic;                     -- mm_interconnect_0:LCD_avalon_slave_read -> LCD:Read_SI
	signal mm_interconnect_0_lcd_avalon_slave_byteenable                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LCD_avalon_slave_byteenable -> LCD:ByteEnable_DI
	signal mm_interconnect_0_lcd_avalon_slave_readdatavalid                    : std_logic;                     -- LCD:ReadDataValid_SO -> mm_interconnect_0:LCD_avalon_slave_readdatavalid
	signal mm_interconnect_0_lcd_avalon_slave_write                            : std_logic;                     -- mm_interconnect_0:LCD_avalon_slave_write -> LCD:Write_SI
	signal mm_interconnect_0_lcd_avalon_slave_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:LCD_avalon_slave_writedata -> LCD:WriteData_DI
	signal mm_interconnect_0_lcd_avalon_slave_burstcount                       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:LCD_avalon_slave_burstcount -> LCD:BurstCount_DI
	signal mm_interconnect_0_sysid_control_slave_readdata                      : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_performance_counter_0_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	signal mm_interconnect_0_performance_counter_0_control_slave_address       : std_logic_vector(4 downto 0);  -- mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	signal mm_interconnect_0_performance_counter_0_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	signal mm_interconnect_0_performance_counter_0_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	signal mm_interconnect_0_performance_counter_0_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                      : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                   : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                   : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                          : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                         : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                       : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                           : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                          : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_altpll_signaltap_pll_slave_readdata               : std_logic_vector(31 downto 0); -- altpll_signalTap:readdata -> mm_interconnect_0:altpll_signalTap_pll_slave_readdata
	signal mm_interconnect_0_altpll_signaltap_pll_slave_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_signalTap_pll_slave_address -> altpll_signalTap:address
	signal mm_interconnect_0_altpll_signaltap_pll_slave_read                   : std_logic;                     -- mm_interconnect_0:altpll_signalTap_pll_slave_read -> altpll_signalTap:read
	signal mm_interconnect_0_altpll_signaltap_pll_slave_write                  : std_logic;                     -- mm_interconnect_0:altpll_signalTap_pll_slave_write -> altpll_signalTap:write
	signal mm_interconnect_0_altpll_signaltap_pll_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_signalTap_pll_slave_writedata -> altpll_signalTap:writedata
	signal mm_interconnect_0_sdram_ctrl_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_chipselect -> SDRAM_ctrl:az_cs
	signal mm_interconnect_0_sdram_ctrl_s1_readdata                            : std_logic_vector(15 downto 0); -- SDRAM_ctrl:za_data -> mm_interconnect_0:SDRAM_ctrl_s1_readdata
	signal mm_interconnect_0_sdram_ctrl_s1_waitrequest                         : std_logic;                     -- SDRAM_ctrl:za_waitrequest -> mm_interconnect_0:SDRAM_ctrl_s1_waitrequest
	signal mm_interconnect_0_sdram_ctrl_s1_address                             : std_logic_vector(22 downto 0); -- mm_interconnect_0:SDRAM_ctrl_s1_address -> SDRAM_ctrl:az_addr
	signal mm_interconnect_0_sdram_ctrl_s1_read                                : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_read -> mm_interconnect_0_sdram_ctrl_s1_read:in
	signal mm_interconnect_0_sdram_ctrl_s1_byteenable                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_ctrl_s1_byteenable -> mm_interconnect_0_sdram_ctrl_s1_byteenable:in
	signal mm_interconnect_0_sdram_ctrl_s1_readdatavalid                       : std_logic;                     -- SDRAM_ctrl:za_valid -> mm_interconnect_0:SDRAM_ctrl_s1_readdatavalid
	signal mm_interconnect_0_sdram_ctrl_s1_write                               : std_logic;                     -- mm_interconnect_0:SDRAM_ctrl_s1_write -> mm_interconnect_0_sdram_ctrl_s1_write:in
	signal mm_interconnect_0_sdram_ctrl_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_ctrl_s1_writedata -> SDRAM_ctrl:az_data
	signal mm_interconnect_0_timer_0_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                               : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                  : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_tcim_s2_chipselect                                : std_logic;                     -- mm_interconnect_0:TCIM_s2_chipselect -> TCIM:chipselect2
	signal mm_interconnect_0_tcim_s2_readdata                                  : std_logic_vector(31 downto 0); -- TCIM:readdata2 -> mm_interconnect_0:TCIM_s2_readdata
	signal mm_interconnect_0_tcim_s2_address                                   : std_logic_vector(9 downto 0);  -- mm_interconnect_0:TCIM_s2_address -> TCIM:address2
	signal mm_interconnect_0_tcim_s2_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:TCIM_s2_byteenable -> TCIM:byteenable2
	signal mm_interconnect_0_tcim_s2_write                                     : std_logic;                     -- mm_interconnect_0:TCIM_s2_write -> TCIM:write2
	signal mm_interconnect_0_tcim_s2_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:TCIM_s2_writedata -> TCIM:writedata2
	signal mm_interconnect_0_tcim_s2_clken                                     : std_logic;                     -- mm_interconnect_0:TCIM_s2_clken -> TCIM:clken2
	signal cpu_tightly_coupled_data_master_0_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_1:CPU_tightly_coupled_data_master_0_readdata -> CPU:dtcm0_readdata
	signal cpu_tightly_coupled_data_master_0_address                           : std_logic_vector(25 downto 0); -- CPU:dtcm0_address -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_address
	signal cpu_tightly_coupled_data_master_0_read                              : std_logic;                     -- CPU:dtcm0_read -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_read
	signal cpu_tightly_coupled_data_master_0_byteenable                        : std_logic_vector(3 downto 0);  -- CPU:dtcm0_byteenable -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_byteenable
	signal cpu_tightly_coupled_data_master_0_write                             : std_logic;                     -- CPU:dtcm0_write -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_write
	signal cpu_tightly_coupled_data_master_0_writedata                         : std_logic_vector(31 downto 0); -- CPU:dtcm0_writedata -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_writedata
	signal cpu_tightly_coupled_data_master_0_clken                             : std_logic;                     -- CPU:dtcm0_clken -> mm_interconnect_1:CPU_tightly_coupled_data_master_0_clken
	signal mm_interconnect_1_tcdm_s1_chipselect                                : std_logic;                     -- mm_interconnect_1:TCDM_s1_chipselect -> TCDM:chipselect
	signal mm_interconnect_1_tcdm_s1_readdata                                  : std_logic_vector(31 downto 0); -- TCDM:readdata -> mm_interconnect_1:TCDM_s1_readdata
	signal mm_interconnect_1_tcdm_s1_address                                   : std_logic_vector(9 downto 0);  -- mm_interconnect_1:TCDM_s1_address -> TCDM:address
	signal mm_interconnect_1_tcdm_s1_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_1:TCDM_s1_byteenable -> TCDM:byteenable
	signal mm_interconnect_1_tcdm_s1_write                                     : std_logic;                     -- mm_interconnect_1:TCDM_s1_write -> TCDM:write
	signal mm_interconnect_1_tcdm_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:TCDM_s1_writedata -> TCDM:writedata
	signal mm_interconnect_1_tcdm_s1_clken                                     : std_logic;                     -- mm_interconnect_1:TCDM_s1_clken -> TCDM:clken
	signal cpu_tightly_coupled_instruction_master_0_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_2:CPU_tightly_coupled_instruction_master_0_readdata -> CPU:itcm0_readdata
	signal cpu_tightly_coupled_instruction_master_0_address                    : std_logic_vector(25 downto 0); -- CPU:itcm0_address -> mm_interconnect_2:CPU_tightly_coupled_instruction_master_0_address
	signal cpu_tightly_coupled_instruction_master_0_read                       : std_logic;                     -- CPU:itcm0_read -> mm_interconnect_2:CPU_tightly_coupled_instruction_master_0_read
	signal cpu_tightly_coupled_instruction_master_0_clken                      : std_logic;                     -- CPU:itcm0_clken -> mm_interconnect_2:CPU_tightly_coupled_instruction_master_0_clken
	signal mm_interconnect_2_tcim_s1_chipselect                                : std_logic;                     -- mm_interconnect_2:TCIM_s1_chipselect -> TCIM:chipselect
	signal mm_interconnect_2_tcim_s1_readdata                                  : std_logic_vector(31 downto 0); -- TCIM:readdata -> mm_interconnect_2:TCIM_s1_readdata
	signal mm_interconnect_2_tcim_s1_address                                   : std_logic_vector(9 downto 0);  -- mm_interconnect_2:TCIM_s1_address -> TCIM:address
	signal mm_interconnect_2_tcim_s1_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_2:TCIM_s1_byteenable -> TCIM:byteenable
	signal mm_interconnect_2_tcim_s1_write                                     : std_logic;                     -- mm_interconnect_2:TCIM_s1_write -> TCIM:write
	signal mm_interconnect_2_tcim_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_2:TCIM_s1_writedata -> TCIM:writedata
	signal mm_interconnect_2_tcim_s1_clken                                     : std_logic;                     -- mm_interconnect_2:TCIM_s1_clken -> TCIM:clken
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [TCDM:reset, TCIM:reset, TCIM:reset2, altpll_signalTap:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, mm_interconnect_1:CPU_reset_reset_bridge_in_reset_reset, mm_interconnect_2:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, TCDM:reset_req, TCIM:reset_req, TCIM:reset_req2, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                       : std_logic;                     -- CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv        : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_ctrl_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_ctrl_s1_read:inv -> SDRAM_ctrl:az_rd_n
	signal mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv                : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_ctrl_s1_byteenable:inv -> SDRAM_ctrl:az_be_n
	signal mm_interconnect_0_sdram_ctrl_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_ctrl_s1_write:inv -> SDRAM_ctrl:az_wr_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, LCD:Reset_NRI, SDRAM_ctrl:reset_n, jtag_uart:rst_n, performance_counter_0:reset_n, sysid:reset_n, timer_0:reset_n]

begin

	cpu : component systemFile_CPU
		port map (
			clk                                 => altpll_0_c0_clk,                                   --                                  clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                                reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                                     .reset_req
			d_address                           => cpu_data_master_address,                           --                          data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                                     .byteenable
			d_read                              => cpu_data_master_read,                              --                                     .read
			d_readdata                          => cpu_data_master_readdata,                          --                                     .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                                     .waitrequest
			d_write                             => cpu_data_master_write,                             --                                     .write
			d_writedata                         => cpu_data_master_writedata,                         --                                     .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                                     .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                                     .debugaccess
			i_address                           => cpu_instruction_master_address,                    --                   instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                                     .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                                     .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                                     .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                                     .readdatavalid
			dtcm0_readdata                      => cpu_tightly_coupled_data_master_0_readdata,        --        tightly_coupled_data_master_0.readdata
			dtcm0_address                       => cpu_tightly_coupled_data_master_0_address,         --                                     .address
			dtcm0_read                          => cpu_tightly_coupled_data_master_0_read,            --                                     .read
			dtcm0_clken                         => cpu_tightly_coupled_data_master_0_clken,           --                                     .clken
			dtcm0_write                         => cpu_tightly_coupled_data_master_0_write,           --                                     .write
			dtcm0_writedata                     => cpu_tightly_coupled_data_master_0_writedata,       --                                     .writedata
			dtcm0_byteenable                    => cpu_tightly_coupled_data_master_0_byteenable,      --                                     .byteenable
			itcm0_readdata                      => cpu_tightly_coupled_instruction_master_0_readdata, -- tightly_coupled_instruction_master_0.readdata
			itcm0_address                       => cpu_tightly_coupled_instruction_master_0_address,  --                                     .address
			itcm0_read                          => cpu_tightly_coupled_instruction_master_0_read,     --                                     .read
			itcm0_clken                         => cpu_tightly_coupled_instruction_master_0_clken,    --                                     .clken
			irq                                 => cpu_irq_irq,                                       --                                  irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --                  debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --                      debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                                     .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                                     .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                                     .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                                     .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                                     .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                                     .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                                     .writedata
			dummy_ci_port                       => open                                               --            custom_instruction_master.readra
		);

	lcd : component LcdDriver
		port map (
			WaitReq_SO            => mm_interconnect_0_lcd_avalon_slave_waitrequest,        -- avalon_slave.waitrequest
			Address_DI            => mm_interconnect_0_lcd_avalon_slave_address,            --             .address
			BurstCount_DI         => mm_interconnect_0_lcd_avalon_slave_burstcount,         --             .burstcount
			ByteEnable_DI         => mm_interconnect_0_lcd_avalon_slave_byteenable,         --             .byteenable
			WriteData_DI          => mm_interconnect_0_lcd_avalon_slave_writedata,          --             .writedata
			ReadData_DO           => mm_interconnect_0_lcd_avalon_slave_readdata,           --             .readdata
			Read_SI               => mm_interconnect_0_lcd_avalon_slave_read,               --             .read
			Write_SI              => mm_interconnect_0_lcd_avalon_slave_write,              --             .write
			ReadDataValid_SO      => mm_interconnect_0_lcd_avalon_slave_readdatavalid,      --             .readdatavalid
			BeginBurstTransfer_SI => mm_interconnect_0_lcd_avalon_slave_beginbursttransfer, --             .beginbursttransfer
			Clk_CI                => altpll_0_c0_clk,                                       --   clock_sink.clk
			Reset_NRI             => rst_controller_reset_out_reset_ports_inv,              --   reset_sink.reset_n
			Cs_NSO                => lcd_conduit_end_cs_n,                                  --  conduit_end.cs_n
			DB_DIO                => lcd_conduit_end_data,                                  --             .data
			DC_NSO                => lcd_conduit_end_data_cmd_n,                            --             .data_cmd_n
			IM0_SO                => lcd_conduit_end_mode,                                  --             .mode
			Rd_NSO                => lcd_conduit_end_rd_n,                                  --             .rd_n
			Wr_NSO                => lcd_conduit_end_wr_n,                                  --             .wr_n
			LcdReset_NRO          => lcd_conduit_end_lcdreset_n                             --             .lcdreset_n
		);

	sdram_ctrl : component systemFile_SDRAM_ctrl
		port map (
			clk            => altpll_0_c0_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,             -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_ctrl_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_ctrl_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_ctrl_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_ctrl_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_ctrl_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_ctrl_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_ctrl_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_ctrl_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_ctrl_wire_addr,                                 --  wire.export
			zs_ba          => sdram_ctrl_wire_ba,                                   --      .export
			zs_cas_n       => sdram_ctrl_wire_cas_n,                                --      .export
			zs_cke         => sdram_ctrl_wire_cke,                                  --      .export
			zs_cs_n        => sdram_ctrl_wire_cs_n,                                 --      .export
			zs_dq          => sdram_ctrl_wire_dq,                                   --      .export
			zs_dqm         => sdram_ctrl_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_ctrl_wire_ras_n,                                --      .export
			zs_we_n        => sdram_ctrl_wire_we_n                                  --      .export
		);

	tcdm : component systemFile_TCDM
		port map (
			clk        => altpll_0_c0_clk,                      --   clk1.clk
			address    => mm_interconnect_1_tcdm_s1_address,    --     s1.address
			clken      => mm_interconnect_1_tcdm_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_tcdm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_tcdm_s1_write,      --       .write
			readdata   => mm_interconnect_1_tcdm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_tcdm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_tcdm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze     => '0'                                   -- (terminated)
		);

	tcim : component systemFile_TCIM
		port map (
			clk         => altpll_0_c0_clk,                      --   clk1.clk
			address     => mm_interconnect_2_tcim_s1_address,    --     s1.address
			clken       => mm_interconnect_2_tcim_s1_clken,      --       .clken
			chipselect  => mm_interconnect_2_tcim_s1_chipselect, --       .chipselect
			write       => mm_interconnect_2_tcim_s1_write,      --       .write
			readdata    => mm_interconnect_2_tcim_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_2_tcim_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_2_tcim_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,   --       .reset_req
			address2    => mm_interconnect_0_tcim_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_tcim_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_tcim_s2_clken,      --       .clken
			write2      => mm_interconnect_0_tcim_s2_write,      --       .write
			readdata2   => mm_interconnect_0_tcim_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_tcim_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_tcim_s2_byteenable, --       .byteenable
			clk2        => altpll_0_c0_clk,                      --   clk2.clk
			reset2      => rst_controller_reset_out_reset,       -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze      => '0'                                   -- (terminated)
		);

	altpll_0 : component systemFile_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,             -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c2                 => altpll_0_c2_clk,                                --                    c2.clk
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			locked             => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "0000",                                         --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	altpll_signaltap : component systemFile_altpll_signalTap
		port map (
			clk                => altpll_0_c0_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                         -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_signaltap_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_signaltap_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_signaltap_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_signaltap_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_signaltap_pll_slave_writedata, --                      .writedata
			c0                 => altpll_1_c0_clk,                                        --                    c0.clk
			scandone           => open,                                                   --           (terminated)
			scandataout        => open,                                                   --           (terminated)
			areset             => '0',                                                    --           (terminated)
			locked             => open,                                                   --           (terminated)
			phasedone          => open,                                                   --           (terminated)
			phasecounterselect => "0000",                                                 --           (terminated)
			phaseupdown        => '0',                                                    --           (terminated)
			phasestep          => '0',                                                    --           (terminated)
			scanclk            => '0',                                                    --           (terminated)
			scanclkena         => '0',                                                    --           (terminated)
			scandata           => '0',                                                    --           (terminated)
			configupdate       => '0'                                                     --           (terminated)
		);

	jtag_uart : component systemFile_jtag_uart
		port map (
			clk            => altpll_0_c0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	performance_counter_0 : component systemFile_performance_counter_0
		port map (
			clk           => altpll_0_c0_clk,                                                     --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                            --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_0_control_slave_writedata      --              .writedata
		);

	sysid : component systemFile_sysid
		port map (
			clock    => altpll_0_c0_clk,                                  --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_0 : component systemFile_timer_0
		port map (
			clk        => altpll_0_c0_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component systemFile_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                            => altpll_0_c0_clk,                                                     --                                          altpll_0_c0.clk
			clk_0_clk_clk                                              => clk_clk,                                                             --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                  -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			CPU_reset_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                                      --                      CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                                    => cpu_data_master_address,                                             --                                      CPU_data_master.address
			CPU_data_master_waitrequest                                => cpu_data_master_waitrequest,                                         --                                                     .waitrequest
			CPU_data_master_byteenable                                 => cpu_data_master_byteenable,                                          --                                                     .byteenable
			CPU_data_master_read                                       => cpu_data_master_read,                                                --                                                     .read
			CPU_data_master_readdata                                   => cpu_data_master_readdata,                                            --                                                     .readdata
			CPU_data_master_readdatavalid                              => cpu_data_master_readdatavalid,                                       --                                                     .readdatavalid
			CPU_data_master_write                                      => cpu_data_master_write,                                               --                                                     .write
			CPU_data_master_writedata                                  => cpu_data_master_writedata,                                           --                                                     .writedata
			CPU_data_master_debugaccess                                => cpu_data_master_debugaccess,                                         --                                                     .debugaccess
			CPU_instruction_master_address                             => cpu_instruction_master_address,                                      --                               CPU_instruction_master.address
			CPU_instruction_master_waitrequest                         => cpu_instruction_master_waitrequest,                                  --                                                     .waitrequest
			CPU_instruction_master_read                                => cpu_instruction_master_read,                                         --                                                     .read
			CPU_instruction_master_readdata                            => cpu_instruction_master_readdata,                                     --                                                     .readdata
			CPU_instruction_master_readdatavalid                       => cpu_instruction_master_readdatavalid,                                --                                                     .readdatavalid
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,                        --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                          --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                           --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,                       --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,                      --                                                     .writedata
			altpll_signalTap_pll_slave_address                         => mm_interconnect_0_altpll_signaltap_pll_slave_address,                --                           altpll_signalTap_pll_slave.address
			altpll_signalTap_pll_slave_write                           => mm_interconnect_0_altpll_signaltap_pll_slave_write,                  --                                                     .write
			altpll_signalTap_pll_slave_read                            => mm_interconnect_0_altpll_signaltap_pll_slave_read,                   --                                                     .read
			altpll_signalTap_pll_slave_readdata                        => mm_interconnect_0_altpll_signaltap_pll_slave_readdata,               --                                                     .readdata
			altpll_signalTap_pll_slave_writedata                       => mm_interconnect_0_altpll_signaltap_pll_slave_writedata,              --                                                     .writedata
			CPU_debug_mem_slave_address                                => mm_interconnect_0_cpu_debug_mem_slave_address,                       --                                  CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                                  => mm_interconnect_0_cpu_debug_mem_slave_write,                         --                                                     .write
			CPU_debug_mem_slave_read                                   => mm_interconnect_0_cpu_debug_mem_slave_read,                          --                                                     .read
			CPU_debug_mem_slave_readdata                               => mm_interconnect_0_cpu_debug_mem_slave_readdata,                      --                                                     .readdata
			CPU_debug_mem_slave_writedata                              => mm_interconnect_0_cpu_debug_mem_slave_writedata,                     --                                                     .writedata
			CPU_debug_mem_slave_byteenable                             => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                    --                                                     .byteenable
			CPU_debug_mem_slave_waitrequest                            => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                   --                                                     .waitrequest
			CPU_debug_mem_slave_debugaccess                            => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                   --                                                     .debugaccess
			jtag_uart_avalon_jtag_slave_address                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,               --                          jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                 --                                                     .write
			jtag_uart_avalon_jtag_slave_read                           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                  --                                                     .read
			jtag_uart_avalon_jtag_slave_readdata                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,              --                                                     .readdata
			jtag_uart_avalon_jtag_slave_writedata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,             --                                                     .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,           --                                                     .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,            --                                                     .chipselect
			LCD_avalon_slave_address                                   => mm_interconnect_0_lcd_avalon_slave_address,                          --                                     LCD_avalon_slave.address
			LCD_avalon_slave_write                                     => mm_interconnect_0_lcd_avalon_slave_write,                            --                                                     .write
			LCD_avalon_slave_read                                      => mm_interconnect_0_lcd_avalon_slave_read,                             --                                                     .read
			LCD_avalon_slave_readdata                                  => mm_interconnect_0_lcd_avalon_slave_readdata,                         --                                                     .readdata
			LCD_avalon_slave_writedata                                 => mm_interconnect_0_lcd_avalon_slave_writedata,                        --                                                     .writedata
			LCD_avalon_slave_beginbursttransfer                        => mm_interconnect_0_lcd_avalon_slave_beginbursttransfer,               --                                                     .beginbursttransfer
			LCD_avalon_slave_burstcount                                => mm_interconnect_0_lcd_avalon_slave_burstcount,                       --                                                     .burstcount
			LCD_avalon_slave_byteenable                                => mm_interconnect_0_lcd_avalon_slave_byteenable,                       --                                                     .byteenable
			LCD_avalon_slave_readdatavalid                             => mm_interconnect_0_lcd_avalon_slave_readdatavalid,                    --                                                     .readdatavalid
			LCD_avalon_slave_waitrequest                               => mm_interconnect_0_lcd_avalon_slave_waitrequest,                      --                                                     .waitrequest
			performance_counter_0_control_slave_address                => mm_interconnect_0_performance_counter_0_control_slave_address,       --                  performance_counter_0_control_slave.address
			performance_counter_0_control_slave_write                  => mm_interconnect_0_performance_counter_0_control_slave_write,         --                                                     .write
			performance_counter_0_control_slave_readdata               => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --                                                     .readdata
			performance_counter_0_control_slave_writedata              => mm_interconnect_0_performance_counter_0_control_slave_writedata,     --                                                     .writedata
			performance_counter_0_control_slave_begintransfer          => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --                                                     .begintransfer
			SDRAM_ctrl_s1_address                                      => mm_interconnect_0_sdram_ctrl_s1_address,                             --                                        SDRAM_ctrl_s1.address
			SDRAM_ctrl_s1_write                                        => mm_interconnect_0_sdram_ctrl_s1_write,                               --                                                     .write
			SDRAM_ctrl_s1_read                                         => mm_interconnect_0_sdram_ctrl_s1_read,                                --                                                     .read
			SDRAM_ctrl_s1_readdata                                     => mm_interconnect_0_sdram_ctrl_s1_readdata,                            --                                                     .readdata
			SDRAM_ctrl_s1_writedata                                    => mm_interconnect_0_sdram_ctrl_s1_writedata,                           --                                                     .writedata
			SDRAM_ctrl_s1_byteenable                                   => mm_interconnect_0_sdram_ctrl_s1_byteenable,                          --                                                     .byteenable
			SDRAM_ctrl_s1_readdatavalid                                => mm_interconnect_0_sdram_ctrl_s1_readdatavalid,                       --                                                     .readdatavalid
			SDRAM_ctrl_s1_waitrequest                                  => mm_interconnect_0_sdram_ctrl_s1_waitrequest,                         --                                                     .waitrequest
			SDRAM_ctrl_s1_chipselect                                   => mm_interconnect_0_sdram_ctrl_s1_chipselect,                          --                                                     .chipselect
			sysid_control_slave_address                                => mm_interconnect_0_sysid_control_slave_address,                       --                                  sysid_control_slave.address
			sysid_control_slave_readdata                               => mm_interconnect_0_sysid_control_slave_readdata,                      --                                                     .readdata
			TCIM_s2_address                                            => mm_interconnect_0_tcim_s2_address,                                   --                                              TCIM_s2.address
			TCIM_s2_write                                              => mm_interconnect_0_tcim_s2_write,                                     --                                                     .write
			TCIM_s2_readdata                                           => mm_interconnect_0_tcim_s2_readdata,                                  --                                                     .readdata
			TCIM_s2_writedata                                          => mm_interconnect_0_tcim_s2_writedata,                                 --                                                     .writedata
			TCIM_s2_byteenable                                         => mm_interconnect_0_tcim_s2_byteenable,                                --                                                     .byteenable
			TCIM_s2_chipselect                                         => mm_interconnect_0_tcim_s2_chipselect,                                --                                                     .chipselect
			TCIM_s2_clken                                              => mm_interconnect_0_tcim_s2_clken,                                     --                                                     .clken
			timer_0_s1_address                                         => mm_interconnect_0_timer_0_s1_address,                                --                                           timer_0_s1.address
			timer_0_s1_write                                           => mm_interconnect_0_timer_0_s1_write,                                  --                                                     .write
			timer_0_s1_readdata                                        => mm_interconnect_0_timer_0_s1_readdata,                               --                                                     .readdata
			timer_0_s1_writedata                                       => mm_interconnect_0_timer_0_s1_writedata,                              --                                                     .writedata
			timer_0_s1_chipselect                                      => mm_interconnect_0_timer_0_s1_chipselect                              --                                                     .chipselect
		);

	mm_interconnect_1 : component systemFile_mm_interconnect_1
		port map (
			altpll_0_c0_clk                              => altpll_0_c0_clk,                              --                       altpll_0_c0.clk
			CPU_reset_reset_bridge_in_reset_reset        => rst_controller_reset_out_reset,               --   CPU_reset_reset_bridge_in_reset.reset
			CPU_tightly_coupled_data_master_0_address    => cpu_tightly_coupled_data_master_0_address,    -- CPU_tightly_coupled_data_master_0.address
			CPU_tightly_coupled_data_master_0_byteenable => cpu_tightly_coupled_data_master_0_byteenable, --                                  .byteenable
			CPU_tightly_coupled_data_master_0_read       => cpu_tightly_coupled_data_master_0_read,       --                                  .read
			CPU_tightly_coupled_data_master_0_readdata   => cpu_tightly_coupled_data_master_0_readdata,   --                                  .readdata
			CPU_tightly_coupled_data_master_0_write      => cpu_tightly_coupled_data_master_0_write,      --                                  .write
			CPU_tightly_coupled_data_master_0_writedata  => cpu_tightly_coupled_data_master_0_writedata,  --                                  .writedata
			CPU_tightly_coupled_data_master_0_clken      => cpu_tightly_coupled_data_master_0_clken,      --                                  .clken
			TCDM_s1_address                              => mm_interconnect_1_tcdm_s1_address,            --                           TCDM_s1.address
			TCDM_s1_write                                => mm_interconnect_1_tcdm_s1_write,              --                                  .write
			TCDM_s1_readdata                             => mm_interconnect_1_tcdm_s1_readdata,           --                                  .readdata
			TCDM_s1_writedata                            => mm_interconnect_1_tcdm_s1_writedata,          --                                  .writedata
			TCDM_s1_byteenable                           => mm_interconnect_1_tcdm_s1_byteenable,         --                                  .byteenable
			TCDM_s1_chipselect                           => mm_interconnect_1_tcdm_s1_chipselect,         --                                  .chipselect
			TCDM_s1_clken                                => mm_interconnect_1_tcdm_s1_clken               --                                  .clken
		);

	mm_interconnect_2 : component systemFile_mm_interconnect_2
		port map (
			altpll_0_c0_clk                                   => altpll_0_c0_clk,                                   --                              altpll_0_c0.clk
			CPU_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                    --          CPU_reset_reset_bridge_in_reset.reset
			CPU_tightly_coupled_instruction_master_0_address  => cpu_tightly_coupled_instruction_master_0_address,  -- CPU_tightly_coupled_instruction_master_0.address
			CPU_tightly_coupled_instruction_master_0_read     => cpu_tightly_coupled_instruction_master_0_read,     --                                         .read
			CPU_tightly_coupled_instruction_master_0_readdata => cpu_tightly_coupled_instruction_master_0_readdata, --                                         .readdata
			CPU_tightly_coupled_instruction_master_0_clken    => cpu_tightly_coupled_instruction_master_0_clken,    --                                         .clken
			TCIM_s1_address                                   => mm_interconnect_2_tcim_s1_address,                 --                                  TCIM_s1.address
			TCIM_s1_write                                     => mm_interconnect_2_tcim_s1_write,                   --                                         .write
			TCIM_s1_readdata                                  => mm_interconnect_2_tcim_s1_readdata,                --                                         .readdata
			TCIM_s1_writedata                                 => mm_interconnect_2_tcim_s1_writedata,               --                                         .writedata
			TCIM_s1_byteenable                                => mm_interconnect_2_tcim_s1_byteenable,              --                                         .byteenable
			TCIM_s1_chipselect                                => mm_interconnect_2_tcim_s1_chipselect,              --                                         .chipselect
			TCIM_s1_clken                                     => mm_interconnect_2_tcim_s1_clken                    --                                         .clken
		);

	irq_mapper : component systemFile_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component systemfile_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => altpll_0_c0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component systemfile_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_ctrl_s1_read_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_read;

	mm_interconnect_0_sdram_ctrl_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_byteenable;

	mm_interconnect_0_sdram_ctrl_s1_write_ports_inv <= not mm_interconnect_0_sdram_ctrl_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of systemFile
